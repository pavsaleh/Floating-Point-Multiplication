--------------------------------------------------------------------------------
-- Title         : 3-bit Adder
-- Project       : VHDL Synthesis Overview
-------------------------------------------------------------------------------
-- File          : threeBitAdder.vhd
-- Author        : Rami Abielmona  <rabielmo@site.uottawa.ca>
-- Created       : 2003/05/17
-- Last modified : 2007/09/25
-------------------------------------------------------------------------------
-- Description : This file creates a 3-bit binary full adder as defined in the VHDL
--		 Synthesis lecture.  The architecture is done at the RTL
--		 abstraction level and the implementation is done in structural
--		 VHDL.
-------------------------------------------------------------------------------
-- Modification history :
-- 2003.05.17 	R. Abielmona		Creation
-- 2004.09.22 	R. Abielmona		Ported for CEG 3550
-- 2007.09.25 	R. Abielmona		Modified copyright notice
-------------------------------------------------------------------------------
-- This file is copyright material of Rami Abielmona, Ph.D., P.Eng., Chief Research
-- Scientist at Larus Technologies.  Permission to make digital or hard copies of part
-- or all of this work for personal or classroom use is granted without fee
-- provided that copies are not made or distributed for profit or commercial
-- advantage and that copies bear this notice and the full citation of this work.
-- Prior permission is required to copy, republish, redistribute or post this work.
-- This notice is adapted from the ACM copyright notice.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY threeBitAdder IS
	PORT (
		i_Ai, i_Bi : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		o_CarryOut : OUT STD_LOGIC;
		o_Sum : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END threeBitAdder;

ARCHITECTURE rtl OF threeBitAdder IS
	SIGNAL int_Sum, int_CarryOut : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL gnd : STD_LOGIC;

	COMPONENT oneBitAdder
		PORT (
			i_CarryIn : IN STD_LOGIC;
			i_Ai, i_Bi : IN STD_LOGIC;
			o_Sum, o_CarryOut : OUT STD_LOGIC);
	END COMPONENT;

BEGIN

	-- Concurrent Signal Assignment
	gnd <= '0';

	add2 : oneBitAdder
	PORT MAP(
		i_CarryIn => gnd,
		i_Ai => i_Ai(2),
		i_Bi => i_Bi(2),
		o_Sum => int_Sum(2),
		o_CarryOut => int_CarryOut(2));

	add1 : oneBitAdder
	PORT MAP(
		i_CarryIn => int_CarryOut(2),
		i_Ai => i_Ai(1),
		i_Bi => i_Bi(1),
		o_Sum => int_Sum(1),
		o_CarryOut => int_CarryOut(1));

	add0 : oneBitAdder
	PORT MAP(
		i_CarryIn => int_CarryOut(1),
		i_Ai => i_Ai(0),
		i_Bi => i_Bi(0),
		o_Sum => int_Sum(0),
		o_CarryOut => int_CarryOut(0));

	-- Output Driver
	o_Sum <= int_Sum;
	o_CarryOut <= int_CarryOut(0);

END rtl;