LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

USE IEEE.STD_LOGIC_ARITH.ALL;

USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY HS IS

    PORT (
        HSA, HSB : IN STD_LOGIC;

        DIFFERENCE, BORROW : OUT STD_LOGIC);

END HS;

ARCHITECTURE dataflow OF HS IS

BEGIN

    DIFFERENCE <= HSA XOR HSB;

    BORROW <= (NOT HSA) AND HSB;

END dataflow;